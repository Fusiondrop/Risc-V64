module ALU #(
    parameter N = 64;
)(
    input   logic [N-1:0] a, b;
    input   logic 
);